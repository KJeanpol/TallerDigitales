module SR_ff_tb();

	reg S_in, R_in, CLK, rst_in;
	wire Q_out;
	
	reg [2:0] testvectors [4:0];
	integer i;

	SR_ff SR_ff_dut(	S_in,
							R_in,
							CLK,
							rst_in,
							Q_out);
							
	initial begin
		$readmemb("C:/Users/kenne/Documents/workspace/Taller Digitales/TallerDigitales/Tarea Flip Flop/JK_ff_testvectors.txt", testvectors);
		i = 0;
	end
	
	always begin
		CLK = 1'b0;
		#5;
		CLK = 1'b1;
		#5;
	end

	always @(posedge CLK) begin
		{S_in, R_in, rst_in} = testvectors[i];
		i = i+1;
	end

endmodule